package apb_tb_pkg;
import uvm_pkg::*;
`include "apb_params.svh"
`include "apb_seq_item.svh"
`include "apb_seqlib.svh"
`include "apb_sequencer.svh"
`include "apb_driver.svh"
`include "apb_monitor.svh"
`include "apb_scoreboard.svh"
`include "apb_agent.svh"
`include "apb_env.svh"
`include "apb_test.svh"
endpackage

`include "apb_checker.sv"
parameter int ADDRESS_WIDTH = 8;
parameter int DATA_WIDTH = 32;